`ifndef STATUS_REGISTER_INDICIES
    `define STATUS_REGISTER_INDICIES 1

    //OPCODE

    `define CARRY_FLAG              0
    `define ZERO_FLAG               1
    `define INTERRUPT_DISABLE_FLAG  2
    `define DECIMAL_MODE_FLAG       3
    `define BRK_FLAG                4
    `define OVERFLOW_FLAG           5
    `define NEGATIVE_FLAG           6
    
`endif
