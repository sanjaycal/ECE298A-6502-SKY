`ifndef REGISTER_IDS

    `define REGISTER_IDS 1
    //OPCODE
    `define ZERO 3'b000
    `define DATA_BUFFER 1
    `define X 2
    `define Y 3
    `define ACC 4
    `define ALU 5
    `define PCH 6
    `define PCL 7

`endif
